-- Copyright (C) 2006 SAMTECH
-- 
-- This library is free software; you can redistribute it and/or
-- modify it under the terms of the GNU Lesser General Public
-- License as published by the Free Software Foundation; either 
-- version 2.1 of the License.
-- 
-- This library is distributed in the hope that it will be useful 
-- but WITHOUT ANY WARRANTY; without even the implied warranty of 
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU 
-- Lesser General Public License for more details.
--
-- You should have received a copy of the GNU Lesser General Public  
-- License along with this library; if not, write to the Free Software 
-- Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307 USA
--
-- See http://www.salome-platform.org/ or email : webmaster.salome@opencascade.com
--  
-- File:	NMTDS_Iterator.cdl
-- Created:	Sun May 07 14:58:16 2006
-- Author:	Peter KURNEV
--		<peter@PREFEX>



class Iterator from NMTDS 

	---Purpose: 

uses 
    ShapeEnum from TopAbs, 
    ShapesDataStructure  from NMTDS,
    PShapesDataStructure from NMTDS,
    ListOfPassKeyBoolean from NMTDS,
    ListIteratorOfListOfPassKeyBoolean from NMTDS
--raises

is 
    Create   
    	returns Iterator from NMTDS;
    ---C++: alias "Standard_EXPORT virtual ~NMTDS_Iterator();" 
    
   
    SetDS(me:out; 
    	    pDS:PShapesDataStructure from NMTDS); 
     
    DS(me) 
      returns ShapesDataStructure from NMTDS; 
    ---C++:return const & 
     
    Initialize(me: out;  
    	    aType1: ShapeEnum from TopAbs;
    	    aType2: ShapeEnum from TopAbs); 
    More(me)  
    	returns Boolean from Standard; 
  	 
    Next(me: out); 
     
    Current(me; aIndex1:out Integer from Standard;
    	    	aIndex2:out Integer from Standard;
    	    	aWithSubShape: out Boolean from Standard); 
    	
    Prepare(me:out); 
     
    ExpectedLength(me) 
    	returns Integer from Standard; 
	 
fields
    myPDS      :PShapesDataStructure from NMTDS     is protected; 
    myLists    :ListOfPassKeyBoolean from NMTDS [6] is protected;  
    myIterator :ListIteratorOfListOfPassKeyBoolean from NMTDS is protected; 
    myEmptyList:ListOfPassKeyBoolean from NMTDS is protected; 
    myLength   :Integer from Standard is protected; 
     
end Iterator;
